module main

import srackham.rimu

fn main() {
	println(rimu.render('*Hello Rimu*!', rimu.RenderOptions{}))
}
